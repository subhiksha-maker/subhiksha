
module Multiplier2x3 (
    input  [1:0] m,
    input  [2:0] q,
    
    output [4:0] p
);


endmodule

